// ---------------------------------------------------------------------------
// File Name :    tb_pkg.svh
// Description :  tb component Class for calculator testbench
// ---------------------------------------------------------------------------

package vip_component_pkg ;
 
  import types_pkg::*;
 `include "stimgen.svh"
 `include "driver.svh"
 `include "monitor.svh"
 `include "reference.svh"
 `include "comparator.svh"
endpackage:vip_component_pkg
// EOF
