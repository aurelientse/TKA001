LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


PACKAGE GCD_DATAPATH_PKG IS


COMPONENT GCD_MUX IS
GENERIC ( DLEN :POSITIVE:=8);
PORT ( 
      a   : IN  STD_LOGIC_VECTOR (DLEN-1 DOWNTO 0);
      b   : IN  STD_LOGIC_VECTOR (DLEN-1 DOWNTO 0);
      s   : IN  STD_LOGIC;
      x   : OUT STD_LOGIC_VECTOR(DLEN-1 DOWNTO 0)
      );
END COMPONENT GCD_MUX;



COMPONENT GCD_REG IS
GENERIC ( DLEN :POSITIVE:=8);
PORT ( 
      clk    : IN  STD_LOGIC;
      rst_n  : IN  STD_LOGIC;
      Load   : IN  STD_LOGIC;
      d      : IN  STD_LOGIC_VECTOR(DLEN-1 DOWNTO 0);
      q      : OUT STD_LOGIC_VECTOR(DLEN-1 DOWNTO 0)
      );
END COMPONENT GCD_REG;

END PACKAGE GCD_DATAPATH_PKG;
