// ---------------------------------------------------------------------------
// File Name :     prog.sv
// Description :   Program for the calculator testbench
// ---------------------------------------------------------------------------

program automatic prog(pins_if pins_vif, output event test_done);
   

   
endprogram

// EOF
